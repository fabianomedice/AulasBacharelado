CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
25 87 998 719
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
25 87 998 719
143654930 0
0
6 Title:
5 Name:
0
0
0
15
14 Logic Display~
6 375 487 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 HLT
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 372 420 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 OUT
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 371 360 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 SUB
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 374 297 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 ADD
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 371 218 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 LDA
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
10 4-In NAND~
219 289 510 0 5 22
0 11 10 9 7 6
0
0 0 112 0
6 74LS20
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
7734 0 0
0
0
9 Inverter~
13 189 210 0 2 22
0 11 13
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
9914 0 0
0
0
9 Inverter~
13 190 236 0 2 22
0 10 12
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
3747 0 0
0
0
9 Inverter~
13 189 260 0 2 22
0 9 14
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 3 0
1 U
3549 0 0
0
0
9 Inverter~
13 190 284 0 2 22
0 7 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 3 0
1 U
7931 0 0
0
0
10 4-In NAND~
219 287 446 0 5 22
0 11 10 9 8 5
0
0 0 112 0
6 74LS20
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
9325 0 0
0
0
10 4-In NAND~
219 286 385 0 5 22
0 13 12 9 8 4
0
0 0 112 0
6 74LS20
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
8903 0 0
0
0
10 4-In NAND~
219 285 326 0 5 22
0 13 12 14 7 3
0
0 0 112 0
6 74LS20
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
3834 0 0
0
0
10 4-In NAND~
219 284 263 0 5 22
0 13 12 14 8 2
0
0 0 112 0
6 74LS20
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 786447
65 0 0 0 2 1 1 0
1 U
3363 0 0
0
0
8 Hex Key~
166 102 175 0 11 12
0 7 9 10 11 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7668 0 0
0
0
29
1 5 2 0 0 8320 0 5 14 0 0 3
371 236
371 263
311 263
1 5 3 0 0 8320 0 4 13 0 0 3
374 315
374 326
312 326
1 5 4 0 0 8320 0 3 12 0 0 3
371 378
371 385
313 385
1 5 5 0 0 8320 0 2 11 0 0 3
372 438
372 446
314 446
1 5 6 0 0 8320 0 1 6 0 0 3
375 505
375 510
316 510
0 4 7 0 0 4224 0 0 6 18 0 3
196 340
196 524
265 524
0 4 8 0 0 8192 0 0 11 15 0 4
219 399
232 399
232 460
263 460
0 3 9 0 0 4096 0 0 6 11 0 3
216 451
216 515
265 515
0 2 10 0 0 4096 0 0 6 12 0 3
225 442
225 506
265 506
0 1 11 0 0 4096 0 0 6 13 0 3
237 433
237 497
265 497
0 3 9 0 0 12288 0 0 11 14 0 4
159 389
160 389
160 451
263 451
0 2 10 0 0 4224 0 0 11 28 0 3
138 236
138 442
263 442
0 1 11 0 0 4224 0 0 11 29 0 3
124 210
124 433
263 433
0 3 9 0 0 4224 0 0 12 27 0 3
159 260
159 390
262 390
0 4 8 0 0 4224 0 0 12 22 0 3
219 284
219 399
262 399
0 2 12 0 0 4096 0 0 12 20 0 3
243 322
243 381
262 381
0 1 13 0 0 8192 0 0 12 21 0 4
246 312
247 312
247 372
262 372
0 4 7 0 0 0 0 0 13 26 0 3
141 284
141 340
261 340
0 3 14 0 0 4224 0 0 13 23 0 3
226 268
226 331
261 331
0 2 12 0 0 4224 0 0 13 24 0 3
231 236
231 322
261 322
0 1 13 0 0 4224 0 0 13 25 0 3
246 210
246 313
261 313
4 2 8 0 0 0 0 14 10 0 0 4
260 277
219 277
219 284
211 284
3 2 14 0 0 0 0 14 9 0 0 4
260 268
226 268
226 260
210 260
2 2 12 0 0 0 0 14 8 0 0 4
260 259
240 259
240 236
211 236
2 1 13 0 0 0 0 7 14 0 0 4
210 210
252 210
252 250
260 250
1 1 7 0 0 0 0 15 10 0 0 3
111 199
111 284
175 284
2 1 9 0 0 0 0 15 9 0 0 3
105 199
105 260
174 260
3 1 10 0 0 0 0 15 8 0 0 3
99 199
99 236
175 236
4 1 11 0 0 0 0 15 7 0 0 3
93 199
93 210
174 210
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
