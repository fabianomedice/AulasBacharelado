CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 9
25 87 998 719
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
25 87 998 719
177209362 0
0
6 Title:
5 Name:
0
0
0
24
7 Ground~
168 175 530 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
2 +V
167 96 429 0 1 3
0 8
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
14 NO PushButton~
191 152 458 0 2 5
0 7 8
0
0 0 4208 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
12 Hex Display~
7 425 518 0 16 19
10 9 10 11 12 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6153 0 0
0
0
10 Buffer 3S~
219 508 444 0 3 22
0 6 7 9
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U3D
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
5394 0 0
0
0
10 Buffer 3S~
219 453 444 0 3 22
0 5 7 10
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U3C
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
7734 0 0
0
0
10 Buffer 3S~
219 401 441 0 3 22
0 4 7 11
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U3B
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
9914 0 0
0
0
10 Buffer 3S~
219 347 441 0 3 22
0 3 7 12
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U3A
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 589827
65 0 0 0 4 1 3 0
1 U
3747 0 0
0
0
7 Pulser~
4 140 353 0 10 12
0 19 20 13 21 0 0 5 5 2
7
0
0 0 4144 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3549 0 0
0
0
12 Hex Display~
7 406 322 0 18 19
10 6 5 4 3 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7931 0 0
0
0
2 +V
167 662 125 0 1 3
0 14
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9325 0 0
0
0
7 Ground~
168 156 226 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8903 0 0
0
0
2 +V
167 183 220 0 1 3
0 16
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3834 0 0
0
0
2 +V
167 88 126 0 1 3
0 18
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3363 0 0
0
0
12 SPST Switch~
165 125 165 0 2 11
0 15 18
0
0 0 4208 0
0
2 S2
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
7668 0 0
0
0
14 NO PushButton~
191 131 275 0 2 5
0 17 2
0
0 0 4208 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4718 0 0
0
0
7 Ground~
168 114 300 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3874 0 0
0
0
6 74112~
219 589 238 0 7 32
0 14 15 4 15 17 22 3
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U2B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 2 2 0
1 U
6671 0 0
0
0
6 74112~
219 492 239 0 7 32
0 14 15 5 15 17 23 4
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U2A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 1 2 0
1 U
3789 0 0
0
0
6 74112~
219 392 237 0 7 32
0 14 15 6 15 17 24 5
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U1B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 2 1 0
1 U
4871 0 0
0
0
6 74112~
219 291 238 0 7 32
0 14 15 13 15 17 25 6
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U1A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 786464
65 0 0 512 2 1 1 0
1 U
3750 0 0
0
0
9 Resistor~
219 175 495 0 3 5
0 2 7 -1
0
0 0 112 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 156 193 0 3 5
0 2 15 -1
0
0 0 112 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 182 253 0 4 5
0 17 16 0 1
0
0 0 112 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
45
1 0 3 0 0 8192 0 8 0 0 8 3
346 427
346 378
397 378
1 0 4 0 0 12288 0 7 0 0 7 4
400 427
400 406
417 406
417 383
1 0 5 0 0 4096 0 6 0 0 6 3
452 430
452 374
428 374
1 0 6 0 0 8192 0 5 0 0 5 3
507 430
507 364
417 364
1 0 6 0 0 16512 0 10 0 0 40 6
415 346
417 346
417 364
332 364
332 206
327 206
2 0 5 0 0 12432 0 10 0 0 39 4
409 346
409 374
429 374
429 212
3 0 4 0 0 12416 0 10 0 0 38 4
403 346
403 383
532 383
532 211
7 4 3 0 0 12416 0 18 10 0 0 5
613 202
623 202
623 389
397 389
397 346
2 0 7 0 0 8192 0 8 0 0 14 3
335 442
317 442
317 466
2 0 7 0 0 0 0 7 0 0 14 3
389 442
383 442
383 466
2 0 7 0 0 0 0 6 0 0 14 3
441 445
425 445
425 466
2 0 7 0 0 0 0 22 0 0 14 2
175 477
175 466
1 1 2 0 0 4224 0 1 22 0 0 2
175 524
175 513
1 2 7 0 0 4224 0 3 5 0 0 4
169 466
489 466
489 445
496 445
1 2 8 0 0 8320 0 2 3 0 0 3
96 438
96 466
135 466
3 1 9 0 0 4224 0 5 4 0 0 4
507 460
507 559
434 559
434 542
3 2 10 0 0 4224 0 6 4 0 0 4
452 460
452 553
428 553
428 542
3 3 11 0 0 4224 0 7 4 0 0 4
400 457
400 556
422 556
422 542
4 3 12 0 0 12416 0 4 8 0 0 4
416 542
416 549
346 549
346 457
3 3 13 0 0 8320 0 21 9 0 0 4
261 211
217 211
217 344
164 344
1 0 14 0 0 4096 0 18 0 0 24 2
589 175
589 142
1 0 14 0 0 4096 0 19 0 0 24 2
492 176
492 142
1 0 14 0 0 0 0 20 0 0 24 2
392 174
392 142
1 1 14 0 0 8320 0 21 11 0 0 4
291 175
291 142
662 142
662 134
1 1 2 0 0 0 0 23 12 0 0 2
156 211
156 220
2 0 15 0 0 4096 0 23 0 0 34 2
156 175
156 165
2 0 15 0 0 4096 0 20 0 0 28 2
368 201
352 201
4 0 15 0 0 8192 0 20 0 0 32 3
368 219
352 219
352 166
4 0 15 0 0 0 0 19 0 0 30 4
468 221
447 221
447 203
448 203
2 0 15 0 0 0 0 19 0 0 32 3
468 203
448 203
448 166
2 0 15 0 0 0 0 18 0 0 32 2
565 202
551 202
0 4 15 0 0 8320 0 0 18 34 0 5
253 165
253 166
551 166
551 220
565 220
2 0 15 0 0 0 0 21 0 0 34 2
267 202
253 202
1 4 15 0 0 0 0 15 21 0 0 4
142 165
253 165
253 220
267 220
1 2 16 0 0 4224 0 13 24 0 0 3
183 229
183 235
182 235
1 0 17 0 0 4096 0 24 0 0 44 2
182 271
182 283
1 2 18 0 0 4224 0 14 15 0 0 3
88 135
88 165
108 165
7 3 4 0 0 0 0 19 18 0 0 5
516 203
516 204
524 204
524 211
559 211
7 3 5 0 0 0 0 20 19 0 0 4
416 201
426 201
426 212
462 212
7 3 6 0 0 0 0 21 20 0 0 4
315 202
327 202
327 210
362 210
5 0 17 0 0 4096 0 21 0 0 44 2
291 250
291 283
5 0 17 0 0 0 0 20 0 0 44 4
392 249
392 278
393 278
393 283
5 0 17 0 0 0 0 19 0 0 44 2
492 251
492 283
5 1 17 0 0 8320 0 18 16 0 0 3
589 250
589 283
148 283
2 1 2 0 0 128 0 16 17 0 0 2
114 283
114 294
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
52 176 132 200
56 180 128 196
9 CONTE(CP)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
55 477 151 501
59 481 147 497
11 ENABLE (EP)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
55 278 103 302
59 282 99 298
5 CLEAR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
