reg6_inst : reg6 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
