CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 8 100 9
0 66 1024 740
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 66 1024 740
177209362 0
0
6 Title:
5 Name:
0
0
0
14
14 Logic Display~
6 99 270 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
6 74112~
219 112 190 0 7 32
0 4 3 5 6 4 7 2
0
0 0 4720 512
7 74LS112
-3 -60 46 -52
3 U3B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 0 2 2 3 0
1 U
4441 0 0
0
0
7 Pulser~
4 878 107 0 10 12
0 16 17 5 18 0 0 5 5 2
8
0
0 0 4656 512
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3618 0 0
0
0
2 +V
167 795 191 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
14 Logic Display~
6 670 271 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 548 270 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 431 269 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 318 270 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 214 270 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
6 74112~
219 668 190 0 7 32
0 4 7 5 2 4 8 12
0
0 0 4720 180
7 74LS112
-3 -60 46 -52
3 U3A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 0 2 1 3 0
1 U
7931 0 0
0
0
6 74112~
219 546 190 0 7 32
0 4 8 5 12 4 13 9
0
0 0 4720 512
7 74LS112
-3 -60 46 -52
3 U2B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 0 2 2 2 0
1 U
9325 0 0
0
0
6 74112~
219 431 190 0 7 32
0 4 9 5 13 4 14 10
0
0 0 4720 512
7 74LS112
-3 -60 46 -52
3 U2A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 0 2 1 2 0
1 U
8903 0 0
0
0
6 74112~
219 319 190 0 7 32
0 4 10 5 14 4 15 11
0
0 0 4720 512
7 74LS112
-3 -60 46 -52
3 U1B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 0 2 2 1 0
1 U
3834 0 0
0
0
6 74112~
219 216 190 0 7 32
0 4 11 5 15 4 6 3
0
0 0 4720 512
7 74LS112
-3 -60 46 -52
3 U1A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -1610612676
65 0 0 0 2 1 1 0
1 U
3363 0 0
0
0
37
1 0 2 0 0 0 0 1 0 0 2 2
99 288
99 288
0 0 2 0 0 4096 0 0 0 10 0 4
63 154
63 296
99 296
99 281
0 1 3 0 0 4224 0 0 9 9 0 4
176 154
176 296
214 296
214 288
1 0 4 0 0 8192 0 2 0 0 20 3
112 127
112 118
216 118
3 0 5 0 0 12288 0 2 0 0 15 4
142 163
159 163
159 99
261 99
4 6 6 0 0 4224 0 2 14 0 0 2
136 172
186 172
5 5 4 0 0 0 0 14 2 0 0 2
216 202
112 202
6 2 7 0 0 12416 0 2 10 0 0 6
82 172
78 172
78 220
706 220
706 172
692 172
2 7 3 0 0 0 0 2 14 0 0 2
136 154
192 154
7 4 2 0 0 12416 0 2 10 0 0 6
88 154
58 154
58 108
706 108
706 154
692 154
3 0 5 0 0 0 0 10 0 0 15 3
698 163
723 163
723 99
3 0 5 0 0 0 0 11 0 0 15 3
576 163
595 163
595 99
3 0 5 0 0 0 0 12 0 0 15 3
461 163
479 163
479 99
3 0 5 0 0 0 0 13 0 0 15 3
349 163
371 163
371 99
3 3 5 0 0 12416 0 14 3 0 0 6
246 163
261 163
261 99
730 99
730 98
854 98
0 0 4 0 0 4096 0 0 0 20 25 3
667 118
776 118
776 199
1 0 4 0 0 0 0 11 0 0 20 2
546 127
546 118
1 0 4 0 0 0 0 12 0 0 20 2
431 127
431 118
1 0 4 0 0 0 0 13 0 0 20 2
319 127
319 118
1 5 4 0 0 8320 0 14 10 0 0 4
216 127
216 118
668 118
668 124
0 1 8 0 0 4224 0 0 5 30 0 4
622 154
622 297
670 297
670 289
0 1 9 0 0 4224 0 0 6 31 0 4
499 154
499 296
548 296
548 288
0 1 10 0 0 4224 0 0 7 32 0 4
393 154
393 295
431 295
431 287
0 1 11 0 0 4224 0 0 8 33 0 4
273 154
273 296
318 296
318 288
1 1 4 0 0 0 0 10 4 0 0 3
668 199
795 199
795 200
5 1 4 0 0 0 0 11 10 0 0 3
546 202
668 202
668 199
5 5 4 0 0 0 0 12 11 0 0 2
431 202
546 202
5 5 4 0 0 0 0 13 12 0 0 2
319 202
431 202
5 5 4 0 0 0 0 14 13 0 0 2
216 202
319 202
2 6 8 0 0 0 0 11 10 0 0 2
570 154
638 154
2 7 9 0 0 0 0 12 11 0 0 2
455 154
522 154
2 7 10 0 0 0 0 13 12 0 0 2
343 154
407 154
2 7 11 0 0 0 0 14 13 0 0 2
240 154
295 154
4 7 12 0 0 4224 0 11 10 0 0 2
570 172
644 172
4 6 13 0 0 4224 0 12 11 0 0 2
455 172
516 172
4 6 14 0 0 4224 0 13 12 0 0 2
343 172
401 172
4 6 15 0 0 4224 0 14 13 0 0 2
240 172
289 172
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
