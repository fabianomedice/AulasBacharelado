CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 0 30 100 9
0 74 804 576
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 74 804 576
177209362 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 815 52 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
9 2-In XOR~
219 772 101 0 3 22
0 2 7 3
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U4D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
4441 0 0
0
0
9 2-In XOR~
219 722 95 0 3 22
0 2 8 4
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U4C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
3618 0 0
0
0
9 2-In XOR~
219 676 91 0 3 22
0 2 9 5
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U4B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
6153 0 0
0
0
9 2-In XOR~
219 626 89 0 3 22
0 2 10 6
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U4A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 571 86 0 3 22
0 2 15 11
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U3D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 527 84 0 3 22
0 2 16 12
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U3C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 486 81 0 3 22
0 2 17 13
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U3B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 439 81 0 3 22
0 2 18 14
0
0 0 112 270
6 74LS86
-21 -24 21 -16
3 U3A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 589837
65 0 0 0 4 1 1 0
1 U
3549 0 0
0
0
14 Logic Display~
6 107 179 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
12 Hex Display~
7 397 251 0 18 19
10 19 20 21 22 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9325 0 0
0
0
12 Hex Display~
7 303 254 0 18 19
10 23 24 25 26 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8903 0 0
0
0
8 Hex Key~
166 683 33 0 11 12
0 7 8 9 10 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3834 0 0
0
0
8 Hex Key~
166 393 30 0 11 12
0 15 16 17 18 0 0 0 0 0
12 67
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3363 0 0
0
0
8 Hex Key~
166 230 53 0 11 12
0 29 30 31 32 0 0 0 0 0
11 66
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7668 0 0
0
0
8 Hex Key~
166 180 53 0 11 12
0 33 34 35 36 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4718 0 0
0
0
6 74LS83
105 475 212 0 14 29
0 32 31 30 29 6 5 4 3 2
22 21 20 19 28
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U2
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
6 74LS83
105 221 190 0 14 29
0 36 35 34 33 14 13 12 11 28
26 25 24 23 27
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U1
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 -1610612668
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
43
9 0 2 0 0 8320 0 17 0 0 2 5
518 182
518 130
761 130
761 74
784 74
1 0 2 0 0 0 0 2 0 0 3 2
784 82
784 47
1 0 2 0 0 0 0 3 0 0 4 3
734 76
734 47
789 47
1 0 2 0 0 0 0 4 0 0 5 4
688 72
688 5
789 5
789 62
1 0 2 0 0 0 0 5 0 0 6 3
638 70
638 62
791 62
1 0 2 0 0 0 0 6 0 0 8 7
583 67
583 55
663 55
663 62
791 62
791 55
796 55
1 0 2 0 0 0 0 7 0 0 8 5
539 65
539 53
663 53
663 62
796 62
1 1 2 0 0 0 0 8 1 0 0 7
498 62
498 52
663 52
663 62
796 62
796 52
801 52
1 1 2 0 0 0 0 9 1 0 0 7
451 62
451 52
663 52
663 62
796 62
796 52
801 52
3 8 3 0 0 8320 0 2 17 0 0 4
775 131
775 174
500 174
500 182
3 7 4 0 0 8320 0 3 17 0 0 4
725 125
725 174
491 174
491 182
3 6 5 0 0 8320 0 4 17 0 0 4
679 121
679 174
482 174
482 182
3 5 6 0 0 8320 0 5 17 0 0 4
629 119
629 174
473 174
473 182
1 2 7 0 0 8320 0 13 2 0 0 4
692 57
692 63
766 63
766 82
2 2 8 0 0 8336 0 13 3 0 0 4
686 57
686 63
716 63
716 76
3 2 9 0 0 8320 0 13 4 0 0 6
680 57
680 62
663 62
663 62
670 62
670 72
4 2 10 0 0 8320 0 13 5 0 0 6
674 57
674 53
614 53
614 57
620 57
620 70
3 8 11 0 0 8320 0 6 18 0 0 4
574 116
574 152
246 152
246 160
3 7 12 0 0 8320 0 7 18 0 0 4
530 114
530 152
237 152
237 160
3 6 13 0 0 8320 0 8 18 0 0 4
489 111
489 152
228 152
228 160
3 5 14 0 0 8320 0 9 18 0 0 4
442 111
442 152
219 152
219 160
1 2 15 0 0 16512 0 14 6 0 0 6
402 54
402 58
430 58
430 51
565 51
565 67
2 2 16 0 0 16512 0 14 7 0 0 6
396 54
396 58
430 58
430 51
521 51
521 65
3 2 17 0 0 16512 0 14 8 0 0 6
390 54
390 58
430 58
430 51
480 51
480 62
4 2 18 0 0 8320 0 14 9 0 0 6
384 54
384 58
430 58
430 51
433 51
433 62
13 1 19 0 0 8320 0 17 11 0 0 4
491 246
491 311
406 311
406 275
12 2 20 0 0 8320 0 17 11 0 0 4
482 246
482 297
400 297
400 275
11 3 21 0 0 8320 0 17 11 0 0 4
473 246
473 291
394 291
394 275
10 4 22 0 0 8320 0 17 11 0 0 4
464 246
464 283
388 283
388 275
13 1 23 0 0 8320 0 18 12 0 0 4
237 224
237 296
312 296
312 278
12 2 24 0 0 8320 0 18 12 0 0 4
228 224
228 286
306 286
306 278
11 3 25 0 0 8320 0 18 12 0 0 3
219 224
219 278
300 278
10 4 26 0 0 8320 0 18 12 0 0 4
210 224
210 272
294 272
294 278
14 1 27 0 0 8320 0 18 10 0 0 6
264 224
264 232
106 232
106 215
107 215
107 197
14 9 28 0 0 8320 0 17 18 0 0 6
518 246
518 213
279 213
279 154
264 154
264 160
1 4 29 0 0 8320 0 15 17 0 0 4
239 77
239 121
464 121
464 182
2 3 30 0 0 8320 0 15 17 0 0 4
233 77
233 129
455 129
455 182
3 2 31 0 0 8320 0 15 17 0 0 4
227 77
227 137
446 137
446 182
4 1 32 0 0 8320 0 15 17 0 0 4
221 77
221 145
437 145
437 182
1 4 33 0 0 12416 0 16 18 0 0 4
189 77
189 103
210 103
210 160
2 3 34 0 0 12416 0 16 18 0 0 4
183 77
183 109
201 109
201 160
3 2 35 0 0 12416 0 16 18 0 0 4
177 77
177 113
192 113
192 160
4 1 36 0 0 12416 0 16 18 0 0 4
171 77
171 117
183 117
183 160
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
