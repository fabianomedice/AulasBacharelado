CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 74 1024 734
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 74 1024 734
177209362 0
0
6 Title:
5 Name:
0
0
0
10
7 Ground~
168 450 133 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
14 Logic Display~
6 107 179 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
12 Hex Display~
7 397 251 0 18 19
10 3 4 5 6 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3618 0 0
0
0
12 Hex Display~
7 303 254 0 16 19
10 7 8 9 10 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6153 0 0
0
0
8 Hex Key~
166 369 58 0 11 12
0 13 14 15 16 0 0 0 0 0
11 66
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5394 0 0
0
0
8 Hex Key~
166 313 56 0 11 12
0 17 18 19 20 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7734 0 0
0
0
8 Hex Key~
166 230 53 0 11 12
0 21 22 23 24 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9914 0 0
0
0
8 Hex Key~
166 180 53 0 11 12
0 25 26 27 28 0 0 0 0 0
10 65
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3747 0 0
0
0
6 74LS83
105 359 156 0 14 29
0 24 23 22 21 16 15 14 13 2
6 5 4 3 12
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U2
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
6 74LS83
105 221 155 0 14 29
0 28 27 26 25 20 19 18 17 12
10 9 8 7 11
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U1
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 -1610612668
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
27
13 1 3 0 0 4224 0 9 3 0 0 4
375 190
375 311
406 311
406 275
12 2 4 0 0 4224 0 9 3 0 0 4
366 190
366 297
400 297
400 275
11 3 5 0 0 4224 0 9 3 0 0 4
357 190
357 291
394 291
394 275
10 4 6 0 0 4224 0 9 3 0 0 4
348 190
348 283
388 283
388 275
13 1 7 0 0 4224 0 10 4 0 0 4
237 189
237 296
312 296
312 278
12 2 8 0 0 4224 0 10 4 0 0 4
228 189
228 286
306 286
306 278
11 3 9 0 0 4224 0 10 4 0 0 3
219 189
219 278
300 278
10 4 10 0 0 8320 0 10 4 0 0 4
210 189
210 272
294 272
294 278
14 1 11 0 0 8320 0 10 2 0 0 6
264 189
264 232
106 232
106 215
107 215
107 197
14 9 12 0 0 8320 0 9 10 0 0 6
402 190
402 213
279 213
279 124
264 124
264 125
1 9 2 0 0 8320 0 1 9 0 0 4
450 127
450 118
402 118
402 126
1 8 13 0 0 4224 0 5 9 0 0 4
378 82
378 118
384 118
384 126
2 7 14 0 0 4224 0 5 9 0 0 4
372 82
372 118
375 118
375 126
3 6 15 0 0 4224 0 5 9 0 0 2
366 82
366 126
4 5 16 0 0 4224 0 5 9 0 0 4
360 82
360 118
357 118
357 126
1 8 17 0 0 8320 0 6 10 0 0 4
322 80
322 117
246 117
246 125
2 7 18 0 0 8320 0 6 10 0 0 4
316 80
316 115
237 115
237 125
3 6 19 0 0 8320 0 6 10 0 0 4
310 80
310 111
228 111
228 125
4 5 20 0 0 8320 0 6 10 0 0 4
304 80
304 109
219 109
219 125
1 4 21 0 0 8320 0 7 9 0 0 4
239 77
239 93
348 93
348 126
2 3 22 0 0 8320 0 7 9 0 0 4
233 77
233 99
339 99
339 126
3 2 23 0 0 8320 0 7 9 0 0 4
227 77
227 104
330 104
330 126
4 1 24 0 0 8320 0 7 9 0 0 4
221 77
221 108
321 108
321 126
1 4 25 0 0 4224 0 8 10 0 0 4
189 77
189 103
210 103
210 125
2 3 26 0 0 4224 0 8 10 0 0 4
183 77
183 109
201 109
201 125
3 2 27 0 0 4224 0 8 10 0 0 4
177 77
177 113
192 113
192 125
4 1 28 0 0 4224 0 8 10 0 0 4
171 77
171 117
183 117
183 125
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
