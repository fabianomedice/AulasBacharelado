CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
20 78 780 559
177209362 0
0
6 Title:
5 Name:
0
0
0
41
2 +V
167 56 501 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 13 485 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
14 NO PushButton~
191 35 448 0 2 5
0 4 2
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3618 0 0
0
0
12 Hex Display~
7 498 475 0 16 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP2
10 -38 45 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6153 0 0
0
0
9 BuffA 3S~
219 588 381 0 3 22
0 9 4 5
0
0 0 112 270
7 74LS125
-24 -51 25 -43
3 U7D
17 -1 38 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 4 7 0
1 U
5394 0 0
0
0
9 BuffA 3S~
219 445 384 0 3 22
0 10 4 6
0
0 0 112 270
7 74LS125
-24 -51 25 -43
3 U7C
17 -1 38 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
7734 0 0
0
0
9 BuffA 3S~
219 291 386 0 3 22
0 11 4 7
0
0 0 112 270
7 74LS125
-24 -51 25 -43
3 U7B
17 -1 38 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
9914 0 0
0
0
9 BuffA 3S~
219 135 387 0 3 22
0 12 4 8
0
0 0 112 270
7 74LS125
-24 -51 25 -43
3 U7A
17 -1 38 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 -1610612720
65 0 0 0 4 1 7 0
1 U
3747 0 0
0
0
7 Ground~
168 17 120 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
2 +V
167 83 15 0 1 3
0 15
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
7 Pulser~
4 699 339 0 10 12
0 37 38 16 39 0 0 5 5 2
7
0
0 0 4656 512
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9325 0 0
0
0
12 Hex Display~
7 351 403 0 18 19
10 9 10 11 12 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8903 0 0
0
0
8 Hex Key~
166 366 31 0 11 12
0 17 18 19 20 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3834 0 0
0
0
9 Inverter~
13 163 76 0 2 22
0 14 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -1610612644
65 0 0 0 6 1 6 0
1 U
3363 0 0
0
0
7 Ground~
168 74 314 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
2 +V
167 13 328 0 1 3
0 23
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
2 +V
167 16 231 0 1 3
0 24
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
7 Ground~
168 75 400 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
14 NO PushButton~
191 41 340 0 2 5
0 21 23
0
0 0 4720 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3789 0 0
0
0
14 NO PushButton~
191 44 241 0 2 5
0 13 24
0
0 0 4720 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4871 0 0
0
0
14 NO PushButton~
191 45 85 0 2 5
0 14 2
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3750 0 0
0
0
5 4013~
219 623 318 0 6 22
0 13 25 16 21 40 9
0
0 0 4208 512
4 4013
10 -60 38 -52
3 U5B
27 -61 48 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 5 0
1 U
8778 0 0
0
0
5 4013~
219 472 320 0 6 22
0 13 26 16 21 41 10
0
0 0 4208 512
4 4013
10 -60 38 -52
3 U5A
27 -61 48 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 5 0
1 U
538 0 0
0
0
5 4013~
219 330 320 0 6 22
0 13 27 16 21 42 11
0
0 0 4208 512
4 4013
10 -60 38 -52
3 U4B
27 -61 48 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 4 0
1 U
6843 0 0
0
0
5 4013~
219 160 323 0 6 22
0 13 28 16 21 43 12
0
0 0 4208 512
4 4013
10 -60 38 -52
3 U4A
27 -61 48 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 -1610612620
65 0 0 512 2 1 4 0
1 U
3136 0 0
0
0
10 2-In NAND~
219 626 201 0 3 22
0 29 30 25
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
5950 0 0
0
0
10 2-In NAND~
219 662 141 0 3 22
0 17 22 29
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
5670 0 0
0
0
10 2-In NAND~
219 586 140 0 3 22
0 14 9 30
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
6828 0 0
0
0
10 2-In NAND~
219 479 202 0 3 22
0 31 32 26
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
6735 0 0
0
0
10 2-In NAND~
219 514 140 0 3 22
0 18 22 31
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U2D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
8365 0 0
0
0
10 2-In NAND~
219 438 139 0 3 22
0 14 10 32
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U2C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
4132 0 0
0
0
10 2-In NAND~
219 294 135 0 3 22
0 14 11 34
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U1D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
4551 0 0
0
0
10 2-In NAND~
219 370 136 0 3 22
0 19 22 33
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U2A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3635 0 0
0
0
10 2-In NAND~
219 336 205 0 3 22
0 33 34 27
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U2B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3973 0 0
0
0
10 2-In NAND~
219 168 197 0 3 22
0 35 36 28
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U1C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
3851 0 0
0
0
10 2-In NAND~
219 201 138 0 3 22
0 20 22 35
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U1B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
8383 0 0
0
0
10 2-In NAND~
219 130 137 0 3 22
0 14 12 36
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U1A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1610612676
65 0 0 0 4 1 1 0
1 U
9334 0 0
0
0
9 Resistor~
219 75 479 0 3 5
0 3 4 1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 83 50 0 4 5
0 14 15 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 76 367 0 3 5
0 2 21 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 74 274 0 3 5
0 2 13 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
69
1 1 3 0 0 4224 0 38 1 0 0 4
75 497
75 518
56 518
56 510
2 0 4 0 0 8192 0 5 0 0 3 5
574 385
574 399
463 399
463 457
372 457
2 0 4 0 0 12416 0 6 0 0 4 4
431 388
372 388
372 457
153 457
2 0 4 0 0 0 0 7 0 0 5 4
277 390
153 390
153 457
88 457
2 0 4 0 0 0 0 8 0 0 6 5
121 391
88 391
88 457
75 457
75 456
1 2 4 0 0 0 0 3 38 0 0 3
52 456
75 456
75 461
2 1 2 0 0 8320 0 3 2 0 0 3
18 456
13 456
13 479
3 1 5 0 0 4224 0 5 4 0 0 4
592 400
592 507
507 507
507 499
3 2 6 0 0 12416 0 6 4 0 0 6
449 403
449 420
529 420
529 519
501 519
501 499
3 3 7 0 0 8320 0 7 4 0 0 4
295 405
295 521
495 521
495 499
4 3 8 0 0 8320 0 4 8 0 0 4
489 499
489 503
139 503
139 406
1 0 9 0 0 8192 0 5 0 0 26 3
592 370
592 366
561 366
1 0 10 0 0 8192 0 6 0 0 27 3
449 373
449 369
417 369
1 0 11 0 0 8192 0 7 0 0 28 3
295 375
295 371
270 371
1 0 12 0 0 8192 0 8 0 0 29 3
139 376
139 372
113 372
1 0 13 0 0 4096 0 24 0 0 42 2
336 263
336 250
2 1 2 0 0 0 0 21 9 0 0 3
28 93
17 93
17 114
0 1 14 0 0 4096 0 0 37 36 0 2
140 93
140 112
0 1 14 0 0 4096 0 0 14 20 0 4
83 77
140 77
140 76
148 76
1 1 14 0 0 0 0 39 21 0 0 3
83 68
83 93
62 93
1 2 15 0 0 4224 0 10 39 0 0 2
83 24
83 32
3 0 16 0 0 4096 0 11 0 0 23 3
675 330
659 330
659 331
3 0 16 0 0 12288 0 22 0 0 24 4
653 300
659 300
659 331
506 331
3 0 16 0 0 0 0 23 0 0 25 4
502 302
506 302
506 331
366 331
3 3 16 0 0 8320 0 25 24 0 0 5
190 305
190 331
368 331
368 302
360 302
1 0 9 0 0 8320 0 12 0 0 58 5
360 427
360 429
561 429
561 288
562 288
2 0 10 0 0 16384 0 12 0 0 59 6
354 427
355 427
355 451
417 451
417 284
418 284
3 0 11 0 0 12288 0 12 0 0 60 5
348 427
348 442
270 442
270 284
269 284
4 0 12 0 0 8320 0 12 0 0 61 5
342 427
342 431
113 431
113 286
111 286
1 1 17 0 0 8320 0 13 27 0 0 4
375 55
375 60
672 60
672 116
2 1 18 0 0 8320 0 13 30 0 0 4
369 55
369 70
524 70
524 115
3 1 19 0 0 8320 0 13 33 0 0 5
363 55
366 55
366 103
380 103
380 111
4 1 20 0 0 8320 0 13 36 0 0 4
357 55
357 85
211 85
211 113
1 0 14 0 0 8192 0 28 0 0 35 3
596 115
596 95
448 95
1 0 14 0 0 0 0 31 0 0 36 4
448 114
448 94
300 94
300 93
1 0 14 0 0 8320 0 32 0 0 19 4
304 110
304 93
140 93
140 77
4 0 21 0 0 8192 0 22 0 0 38 3
629 324
629 340
478 340
4 0 21 0 0 0 0 23 0 0 39 4
478 326
478 340
336 340
336 341
4 0 21 0 0 8320 0 24 0 0 40 3
336 326
336 341
166 341
4 2 21 0 0 0 0 25 40 0 0 4
166 329
166 341
76 341
76 349
1 0 13 0 0 8192 0 22 0 0 42 3
629 261
629 250
478 250
1 0 13 0 0 8320 0 23 0 0 43 3
478 263
478 250
166 250
1 0 13 0 0 0 0 25 0 0 53 4
166 266
166 250
74 250
74 249
2 0 22 0 0 8192 0 27 0 0 45 3
654 116
654 79
506 79
2 0 22 0 0 0 0 30 0 0 46 3
506 115
506 79
362 79
2 0 22 0 0 8320 0 33 0 0 47 4
362 111
362 77
193 77
193 76
2 2 22 0 0 0 0 14 36 0 0 3
184 76
193 76
193 113
1 1 2 0 0 0 0 18 40 0 0 3
75 394
75 385
76 385
1 1 2 0 0 0 0 15 41 0 0 2
74 308
74 292
1 2 23 0 0 4224 0 16 19 0 0 3
13 337
13 348
24 348
1 2 24 0 0 8320 0 17 20 0 0 3
16 240
16 249
27 249
2 1 21 0 0 0 0 40 19 0 0 3
76 349
76 348
58 348
1 2 13 0 0 0 0 20 41 0 0 3
61 249
74 249
74 256
3 2 25 0 0 12416 0 26 22 0 0 5
627 227
627 240
662 240
662 282
653 282
3 2 26 0 0 12416 0 29 23 0 0 5
480 228
480 241
512 241
512 284
502 284
3 2 27 0 0 12416 0 34 24 0 0 5
337 231
337 239
368 239
368 284
360 284
3 2 28 0 0 12416 0 35 25 0 0 5
169 223
169 239
197 239
197 287
190 287
2 6 9 0 0 0 0 28 22 0 0 7
578 115
578 111
562 111
562 288
562 288
562 282
605 282
2 6 10 0 0 12416 0 31 23 0 0 5
430 114
430 110
418 110
418 284
454 284
2 6 11 0 0 12416 0 32 24 0 0 5
286 110
286 106
269 106
269 284
312 284
2 6 12 0 0 0 0 37 25 0 0 5
122 112
122 108
111 108
111 287
142 287
3 1 29 0 0 8320 0 27 26 0 0 4
663 167
663 177
636 177
636 176
3 2 30 0 0 8320 0 28 26 0 0 4
587 166
587 177
618 177
618 176
3 1 31 0 0 8320 0 30 29 0 0 4
515 166
515 176
489 176
489 177
3 2 32 0 0 8320 0 31 29 0 0 4
439 165
439 176
471 176
471 177
3 1 33 0 0 8320 0 33 34 0 0 4
371 162
371 172
346 172
346 180
3 2 34 0 0 8320 0 32 34 0 0 4
295 161
295 172
328 172
328 180
3 1 35 0 0 8320 0 36 35 0 0 4
202 164
202 178
178 178
178 172
2 3 36 0 0 8320 0 35 37 0 0 4
160 172
160 171
131 171
131 163
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
