CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 100 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
20 78 780 559
177209362 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 299 376 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 301 189 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 31 448 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 107 216 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 123 137 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 126 43 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
9 2-In NOR~
219 225 428 0 3 22
0 6 5 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1610612639
65 0 0 0 4 1 5 0
1 U
9914 0 0
0
0
9 Inverter~
13 100 455 0 2 22
0 6 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 -1610612720
65 0 0 0 6 3 2 0
1 U
3747 0 0
0
0
9 2-In AND~
219 177 456 0 3 22
0 8 8 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1610612636
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
9 Inverter~
13 126 288 0 2 22
0 10 9
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
7931 0 0
0
0
10 2-In NAND~
219 191 321 0 3 22
0 7 9 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 189 218 0 3 22
0 10 7 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -1610612636
65 0 0 0 4 3 1 0
1 U
8903 0 0
0
0
14 Logic Display~
6 465 313 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 454 234 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
10 3-In NAND~
219 338 331 0 4 22
0 14 11 3 13
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 3 0
1 U
7668 0 0
0
0
10 3-In NAND~
219 338 255 0 4 22
0 4 12 13 14
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 -1610612628
65 0 0 0 3 1 3 0
1 U
4718 0 0
0
0
7 Ground~
168 421 191 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
9 DC Motor~
219 375 129 0 2 5
0 15 2
0
0 0 624 0
4 100H
-15 -42 13 -34
2 M1
-7 -26 7 -18
0
0
27 %D %1 N%D %V
R%D N%D %2 10
0
0
4 SIP2
5

0 1 2 1 2 -1610612720
76 0 0 0 1 0 0 0
1 M
6671 0 0
0
0
9 Inverter~
13 178 42 0 2 22
0 17 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -1610612720
65 0 0 0 6 1 2 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 256 126 0 3 22
0 19 16 15
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
4871 0 0
0
0
10 2-In NAND~
219 256 58 0 3 22
0 18 15 19
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-15 -43 6 -35
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1610612676
65 0 0 0 4 1 1 0
1 U
3750 0 0
0
0
28
3 1 3 0 0 8320 0 15 1 0 0 6
314 340
310 340
310 366
317 366
317 376
311 376
1 1 4 0 0 8320 0 2 16 0 0 6
313 189
318 189
318 236
309 236
309 246
314 246
2 0 5 0 0 4096 0 7 0 0 8 2
212 437
212 438
1 0 6 0 0 4096 0 7 0 0 5 2
212 419
212 420
0 0 6 0 0 4224 0 0 0 0 6 3
220 420
68 420
68 448
1 1 6 0 0 0 0 3 8 0 0 4
43 448
77 448
77 455
85 455
3 0 7 0 0 12416 0 7 0 0 13 6
264 428
265 428
265 368
89 368
89 273
159 273
0 3 5 0 0 8320 0 0 9 0 0 4
220 438
206 438
206 456
198 456
2 0 8 0 0 4096 0 9 0 0 10 3
153 465
137 465
137 455
2 1 8 0 0 4224 0 8 9 0 0 4
121 455
145 455
145 447
153 447
2 0 9 0 0 4096 0 10 0 0 14 2
129 306
130 330
0 1 10 0 0 4224 0 0 10 15 0 4
130 216
130 262
129 262
129 270
2 1 7 0 0 0 0 12 11 0 0 4
165 227
159 227
159 312
167 312
2 0 9 0 0 4224 0 11 0 0 0 4
167 330
130 330
130 331
121 331
1 1 10 0 0 0 0 4 12 0 0 4
119 216
157 216
157 209
165 209
3 2 11 0 0 4224 0 11 15 0 0 4
218 321
306 321
306 331
314 331
3 2 12 0 0 4224 0 12 16 0 0 4
216 218
306 218
306 255
314 255
1 0 13 0 0 8320 0 13 0 0 20 4
465 331
465 336
378 336
378 331
1 0 14 0 0 8320 0 14 0 0 21 3
454 252
454 258
369 258
4 3 13 0 0 0 0 15 16 0 0 6
365 331
378 331
378 288
306 288
306 264
314 264
4 1 14 0 0 0 0 16 15 0 0 6
365 255
369 255
369 306
306 306
306 322
314 322
1 0 15 0 0 4224 0 18 0 0 27 3
351 128
287 128
287 126
2 1 2 0 0 8320 0 18 17 0 0 3
399 128
421 128
421 185
1 2 16 0 0 4224 0 5 20 0 0 4
135 137
224 137
224 135
232 135
1 1 17 0 0 4224 0 19 6 0 0 4
163 42
147 42
147 43
138 43
2 1 18 0 0 4224 0 19 21 0 0 4
199 42
224 42
224 49
232 49
3 2 15 0 0 0 0 20 21 0 0 6
283 126
287 126
287 78
224 78
224 67
232 67
3 1 19 0 0 12416 0 21 20 0 0 6
283 58
300 58
300 94
224 94
224 117
232 117
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
