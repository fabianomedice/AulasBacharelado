CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
16 72 624 445
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
16 72 624 445
177209362 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 105 254 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
12 Hex Display~
7 319 120 0 18 19
10 2 3 4 5 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4441 0 0
0
0
9 2-In XOR~
219 197 222 0 3 22
0 10 6 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3618 0 0
0
0
9 2-In XOR~
219 194 175 0 3 22
0 9 6 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
6153 0 0
0
0
9 2-In XOR~
219 199 131 0 3 22
0 8 6 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 199 77 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1610612672
65 0 0 0 4 1 1 0
1 U
7734 0 0
0
0
8 Hex Key~
166 104 51 0 11 12
0 7 8 9 10 0 0 0 0 0
11 66
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9914 0 0
0
0
12
1 3 2 0 0 12416 0 2 6 0 0 5
328 144
328 159
248 159
248 77
232 77
2 3 3 0 0 8320 0 2 5 0 0 5
322 144
322 153
240 153
240 131
232 131
3 3 4 0 0 8320 0 2 4 0 0 3
316 144
316 175
227 175
4 3 5 0 0 8320 0 2 3 0 0 3
310 144
310 222
230 222
2 0 6 0 0 4096 0 3 0 0 8 2
181 231
126 231
2 0 6 0 0 0 0 4 0 0 8 2
178 184
126 184
2 0 6 0 0 4096 0 5 0 0 8 2
183 140
126 140
2 1 6 0 0 8320 0 6 1 0 0 4
183 86
126 86
126 254
117 254
1 1 7 0 0 8320 0 7 6 0 0 5
113 75
113 79
175 79
175 68
183 68
2 1 8 0 0 8320 0 7 5 0 0 3
107 75
107 122
183 122
3 1 9 0 0 4224 0 7 4 0 0 3
101 75
101 166
178 166
4 1 10 0 0 4224 0 7 3 0 0 3
95 75
95 213
181 213
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
