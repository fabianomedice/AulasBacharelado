CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 9
25 87 998 719
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
25 87 998 719
177209362 0
0
6 Title:
5 Name:
0
0
0
39
7 Ground~
168 134 670 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
2 +V
167 78 575 0 1 3
0 4
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
14 NO PushButton~
191 109 598 0 2 5
0 3 4
0
0 0 4208 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
12 Hex Display~
7 523 662 0 16 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6153 0 0
0
0
10 Buffer 3S~
219 703 566 0 3 22
0 9 3 5
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U7D
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 4 7 0
1 U
5394 0 0
0
0
10 Buffer 3S~
219 580 565 0 3 22
0 10 3 6
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U7C
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
7734 0 0
0
0
10 Buffer 3S~
219 462 564 0 3 22
0 11 3 7
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U7B
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
9914 0 0
0
0
10 Buffer 3S~
219 310 562 0 3 22
0 12 3 8
0
0 0 112 270
7 74LS126
-24 -51 25 -43
3 U7A
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 589837
65 0 0 0 4 1 7 0
1 U
3747 0 0
0
0
7 Pulser~
4 120 457 0 10 12
0 39 40 13 41 0 0 5 5 1
8
0
0 0 4144 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3549 0 0
0
0
12 Hex Display~
7 516 485 0 18 19
10 9 10 11 12 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7931 0 0
0
0
2 +V
167 858 415 0 1 3
0 14
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9325 0 0
0
0
8 Hex Key~
166 419 59 0 11 12
0 15 16 17 18 0 0 0 0 0
10 65
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
8903 0 0
0
0
10 2-In NAND~
219 220 243 0 3 22
0 12 19 37
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
3834 0 0
0
0
10 2-In NAND~
219 156 245 0 3 22
0 18 20 36
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3363 0 0
0
0
10 2-In NAND~
219 190 303 0 3 22
0 37 36 35
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
7668 0 0
0
0
9 Inverter~
13 182 388 0 2 22
0 35 38
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
4718 0 0
0
0
6 74112~
219 251 406 0 7 32
0 25 35 13 38 14 42 12
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U1A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 1 1 0
1 U
3874 0 0
0
0
6 74112~
219 428 406 0 7 32
0 25 22 13 34 14 43 11
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U1B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 2 1 0
1 U
6671 0 0
0
0
9 Inverter~
13 359 388 0 2 22
0 22 34
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 363 301 0 3 22
0 33 32 22
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U4B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
4871 0 0
0
0
10 2-In NAND~
219 333 244 0 3 22
0 17 20 32
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U4A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 4 0
1 U
3750 0 0
0
0
10 2-In NAND~
219 396 246 0 3 22
0 11 19 33
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U3D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
8778 0 0
0
0
6 74112~
219 611 410 0 7 32
0 25 23 13 31 14 44 10
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U6A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 1 6 0
1 U
538 0 0
0
0
9 Inverter~
13 542 392 0 2 22
0 23 31
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 2 0
1 U
6843 0 0
0
0
10 2-In NAND~
219 544 303 0 3 22
0 30 29 23
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U5A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
3136 0 0
0
0
10 2-In NAND~
219 514 241 0 3 22
0 16 20 29
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U4D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 4 0
1 U
5950 0 0
0
0
10 2-In NAND~
219 573 242 0 3 22
0 10 19 30
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U4C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
5670 0 0
0
0
6 74112~
219 782 410 0 7 32
0 25 24 13 28 14 45 9
0
0 0 4208 0
7 74LS76A
-3 -60 46 -52
3 U6B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 2 6 0
1 U
6828 0 0
0
0
9 Inverter~
13 713 392 0 2 22
0 24 28
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 2 0
1 U
6735 0 0
0
0
10 2-In NAND~
219 714 302 0 3 22
0 27 26 24
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U5D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 5 0
1 U
8365 0 0
0
0
10 2-In NAND~
219 684 244 0 3 22
0 15 20 26
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U5C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 5 0
1 U
4132 0 0
0
0
10 2-In NAND~
219 743 244 0 3 22
0 9 19 27
0
0 0 112 270
6 74LS00
-14 -24 28 -16
3 U5B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
4551 0 0
0
0
2 +V
167 861 300 0 1 3
0 25
0
0 0 53744 0
2 5V
-6 -23 8 -15
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3635 0 0
0
0
14 NO PushButton~
191 79 185 0 2 5
0 20 21
0
0 0 4208 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3973 0 0
0
0
7 Ground~
168 106 253 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3851 0 0
0
0
2 +V
167 53 157 0 1 3
0 21
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8383 0 0
0
0
9 Inverter~
13 138 154 0 2 22
0 20 19
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 2 0
1 U
9334 0 0
0
0
9 Resistor~
219 134 639 0 3 5
0 2 3 -1
0
0 0 112 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 106 222 0 3 5
0 2 20 -1
0
0 0 112 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
71
2 0 3 0 0 4096 0 38 0 0 5 2
134 621
134 606
2 0 3 0 0 4096 0 6 0 0 4 3
568 566
522 566
522 607
2 0 3 0 0 0 0 7 0 0 4 3
450 565
412 565
412 607
0 2 3 0 0 8336 0 0 5 5 0 5
291 606
291 607
684 607
684 567
691 567
1 2 3 0 0 0 0 3 8 0 0 4
126 606
291 606
291 563
298 563
1 1 2 0 0 4224 0 1 38 0 0 2
134 664
134 657
1 2 4 0 0 4224 0 2 3 0 0 3
78 584
78 606
92 606
3 1 5 0 0 8320 0 5 4 0 0 4
702 582
702 694
532 694
532 686
3 2 6 0 0 4224 0 6 4 0 0 4
579 581
579 714
526 714
526 686
3 3 7 0 0 4224 0 7 4 0 0 4
461 580
461 712
520 712
520 686
3 4 8 0 0 8320 0 8 4 0 0 4
309 578
309 694
514 694
514 686
1 0 9 0 0 4096 0 5 0 0 16 2
702 552
702 513
1 0 10 0 0 4096 0 6 0 0 17 2
579 551
579 531
1 0 11 0 0 12288 0 7 0 0 22 4
461 550
461 552
462 552
462 530
1 0 12 0 0 4096 0 8 0 0 23 2
309 548
309 516
1 0 9 0 0 8320 0 10 0 0 51 4
525 509
525 513
825 513
825 370
2 0 10 0 0 12416 0 10 0 0 56 4
519 509
519 531
651 531
651 374
3 0 13 0 0 8192 0 17 0 0 21 3
221 379
217 379
217 448
3 0 13 0 0 0 0 18 0 0 21 3
398 379
390 379
390 448
3 0 13 0 0 0 0 23 0 0 21 3
581 383
567 383
567 448
3 3 13 0 0 4224 0 9 28 0 0 4
144 448
744 448
744 383
752 383
0 3 11 0 0 4224 0 0 10 61 0 4
462 370
462 530
513 530
513 509
4 0 12 0 0 8320 0 10 0 0 66 4
507 509
507 516
285 516
285 370
5 0 14 0 0 4096 0 28 0 0 27 3
782 422
782 432
781 432
5 0 14 0 0 0 0 23 0 0 27 3
611 422
611 432
610 432
5 0 14 0 0 4096 0 18 0 0 27 2
428 418
428 432
5 1 14 0 0 8320 0 17 11 0 0 4
251 418
251 432
858 432
858 424
1 1 15 0 0 8320 0 12 31 0 0 4
428 83
428 106
694 106
694 219
2 1 16 0 0 8320 0 12 26 0 0 4
422 83
422 134
524 134
524 216
3 1 17 0 0 12416 0 12 21 0 0 4
416 83
416 134
343 134
343 219
4 1 18 0 0 8320 0 12 14 0 0 4
410 83
410 108
166 108
166 220
2 0 19 0 0 4096 0 13 0 0 35 2
212 218
212 154
2 0 19 0 0 4096 0 22 0 0 35 2
388 221
388 154
2 0 19 0 0 0 0 27 0 0 35 2
565 217
565 154
2 2 19 0 0 4224 0 37 32 0 0 3
159 154
735 154
735 219
1 0 20 0 0 8192 0 37 0 0 37 4
123 154
107 154
107 193
106 193
2 0 20 0 0 0 0 39 0 0 41 2
106 204
106 193
2 0 20 0 0 0 0 14 0 0 41 2
148 220
148 193
2 0 20 0 0 0 0 21 0 0 41 4
325 219
325 198
326 198
326 193
2 0 20 0 0 0 0 26 0 0 41 2
506 216
506 193
1 2 20 0 0 4224 0 34 31 0 0 3
96 193
676 193
676 219
1 2 21 0 0 4224 0 36 34 0 0 3
53 166
53 193
62 193
1 1 2 0 0 128 0 35 39 0 0 2
106 247
106 240
3 0 22 0 0 4096 0 20 0 0 65 2
364 327
364 370
3 0 23 0 0 4096 0 25 0 0 60 2
545 329
545 374
3 0 24 0 0 4096 0 30 0 0 55 2
715 328
715 374
1 0 25 0 0 4096 0 23 0 0 50 2
611 347
611 333
1 0 25 0 0 0 0 28 0 0 50 2
782 347
782 333
1 0 25 0 0 0 0 18 0 0 50 2
428 343
428 333
1 1 25 0 0 8320 0 17 33 0 0 4
251 343
251 333
861 333
861 309
7 1 9 0 0 0 0 28 32 0 0 5
806 374
825 374
825 215
753 215
753 219
3 2 26 0 0 8320 0 31 30 0 0 3
685 270
685 277
706 277
3 1 27 0 0 8320 0 32 30 0 0 3
744 270
744 277
724 277
2 4 28 0 0 4224 0 29 28 0 0 2
734 392
758 392
2 1 24 0 0 4224 0 28 29 0 0 4
758 374
690 374
690 392
698 392
7 1 10 0 0 8320 0 23 27 0 0 5
635 374
652 374
652 210
583 210
583 217
3 2 29 0 0 8320 0 26 25 0 0 3
515 267
515 278
536 278
3 1 30 0 0 8320 0 27 25 0 0 3
574 268
574 278
554 278
2 4 31 0 0 4224 0 24 23 0 0 2
563 392
587 392
2 1 23 0 0 4224 0 23 24 0 0 4
587 374
519 374
519 392
527 392
7 1 11 0 0 0 0 18 22 0 0 5
452 370
462 370
462 215
406 215
406 221
3 2 32 0 0 8320 0 21 20 0 0 3
334 270
334 276
355 276
3 1 33 0 0 8320 0 22 20 0 0 3
397 272
397 276
373 276
2 4 34 0 0 4224 0 19 18 0 0 2
380 388
404 388
2 1 22 0 0 4224 0 18 19 0 0 4
404 370
336 370
336 388
344 388
7 1 12 0 0 0 0 17 13 0 0 4
275 370
285 370
285 218
230 218
3 0 35 0 0 4096 0 15 0 0 71 2
191 329
191 370
3 2 36 0 0 8320 0 14 15 0 0 3
157 271
157 278
182 278
3 1 37 0 0 8320 0 13 15 0 0 3
221 269
221 278
200 278
2 4 38 0 0 4224 0 16 17 0 0 2
203 388
227 388
2 1 35 0 0 4224 0 17 16 0 0 4
227 370
159 370
159 388
167 388
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
200 570 216 594
204 574 212 590
1 '
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
21 206 93 230
25 210 89 226
8 LOAD (L)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
22 618 110 642
26 622 106 638
10 ENABLE (E)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
